`timescale 1ns/1ns

module song_loader(song_select, output_red, output_blue, output_yellow, output_total_notes);
  input [4:0] song_select;
  output [99:0] output_red, output_blue, output_yellow;
  
  output [7:0] output_total_notes;
  reg [7:0] total_notes;
  assign output_total_notes = total_notes;

  localparam Take_on_Me = 5'b00011, // Songs available
             Through_The_Fire_and_Flames = 5'b11111;
  
  reg [99:0] red, blue, yellow;
  
  assign output_red = red;
  assign output_blue = blue;
  assign output_yellow = yellow;
  
  always @(*)
  begin
    case (song_select[4:0])
      // More cases to be added in future, each case is its own song
      Through_The_Fire_and_Flames:
        begin
          red    <= 100'b0000000000101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010;
          yellow <= 100'b0000000000010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001;
          blue   <= 100'b0000000000000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100;
          total_notes <= 8'd90;
        end
      Take_on_Me:
        begin
          red    <= 100'b0000000000000000000001010101010101010000000000000000010101010000000000000000010101010000000000000000;
          yellow <= 100'b0000000000111111111100000000000000000101010001010101000000000101000001010101000000000000000000000000;
          blue   <= 100'b0000000000011111111100000000000000000000000100000000000000000000010100000000000000000000000000000000;
          total_notes <= 8'd42;
        end
      default:
        begin // Default is no song
          red    <= 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
          yellow <= 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
          blue   <= 100'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
          total_notes <= 0;
        end
    endcase
  end
endmodule
